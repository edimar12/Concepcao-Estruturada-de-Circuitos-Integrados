library verilog;
use verilog.vl_types.all;
entity extend_tb is
end extend_tb;
