library verilog;
use verilog.vl_types.all;
entity inv_tb is
end inv_tb;
