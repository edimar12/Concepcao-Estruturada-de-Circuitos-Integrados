library verilog;
use verilog.vl_types.all;
entity acc_tb is
end acc_tb;
