module mux2(a, b, s, y);
	input logic [3:0] a, b;
	output logic [3:0] y;
	input logic s;
	assign y = s ? b : a;
endmodule