library verilog;
use verilog.vl_types.all;
entity reg_tb is
end reg_tb;
