library verilog;
use verilog.vl_types.all;
entity addacc_tb is
end addacc_tb;
